module tt_franc_simple_inverter(
input wire in,
output wire out);


assign out = ~in;


endmodule
